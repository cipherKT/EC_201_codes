module andgate_tb;
reg a,b;
wire y,p;

andgate uut(y,a,b);

initial begin 
$dumpfile("test_and.vcd");
$dumpvars(0,andgate_tb);


a = 0;
b = 0;
#5
a = 0;
b = 1;
#5
a = 1;
b = 0;
#5
a = 1;
b = 1;
#5
a = 0;
b = 0;
#5
$finish();
end
endmodule

