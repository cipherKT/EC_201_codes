module nandgate(a,b,y);
input a,b;
output y;

nand(y,a,b);

endmodule

