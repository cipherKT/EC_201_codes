module norgate(a,b,y);
input a,b;
output y;
nor(y,a,b);
endmodule
