module notgate_(a,y);
input a;
output y;

not(y,a);

endmodule

