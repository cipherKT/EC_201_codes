module xorgate(a,b,y);
input a,b;
output y;
xor(y,a,b);
endmodule
