module notgate(y,a);
input a;
output y;

nand(y,a,a);

endmodule

